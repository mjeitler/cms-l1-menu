-- ========================================================
-- from VHDL producer:

-- Module ID: 4

-- Name of L1 Trigger Menu:
-- L1Menu_Collisions2018_v2_0_0

-- Unique ID of L1 Trigger Menu:
-- 669da877-bfe2-4b02-842e-13ee40f3e064

-- Unique ID of firmware implementation:
-- cfa03eba-c8d7-4d4f-9e2c-8039338ad141

-- Scale set:
-- scales_2017_05_23

-- VHDL producer version
-- v2.4.0

-- HB 2016-09-16: constants for algo_mapping_rop.
type global_index_array is array (0 to NR_ALGOS-1) of integer;
constant global_index: global_index_array := (
        143, -- module_index: 0, name: L1_DoubleMu3_dR_Max1p6_Jet90er2p5_dR_Max0p8
        126, -- module_index: 1, name: L1_Mu3_Jet120er2p5_dR_Max0p4
        122, -- module_index: 2, name: L1_Mu3_Jet35er2p5_dR_Max0p4
        258, -- module_index: 3, name: L1_LooseIsoEG24er2p1_IsoTau27er2p1_dR_Min0p3
        348, -- module_index: 4, name: L1_DoubleJet30er2p5_Mass_Min150_dEta_Max1p5
        352, -- module_index: 5, name: L1_DoubleJet30er2p5_Mass_Min330_dEta_Max1p5
        359, -- module_index: 6, name: L1_DoubleJet_120_45_DoubleJet45_Mass_Min620
        382, -- module_index: 7, name: L1_QuadJet60er2p5
        494, -- module_index: 8, name: L1_CDC_SingleMu_3_er1p2_TOP120_DPHI2p618_3p142
         59, -- module_index: 9, name: L1_DoubleMu0er1p4_SQ_OS_dR_Max1p4
         61, -- module_index: 10, name: L1_DoubleMu4_SQ_OS_dR_Max1p2
         80, -- module_index: 11, name: L1_TripleMu_5_5_3
         56, -- module_index: 12, name: L1_DoubleMu0er1p5_SQ_OS
         44, -- module_index: 13, name: L1_DoubleMu8_SQ
        104, -- module_index: 14, name: L1_Mu6_DoubleEG10er2p5
        131, -- module_index: 15, name: L1_Mu6_HTT240er
        107, -- module_index: 16, name: L1_Mu6_DoubleEG17er2p5
        106, -- module_index: 17, name: L1_Mu6_DoubleEG15er2p5
        105, -- module_index: 18, name: L1_Mu6_DoubleEG12er2p5
        132, -- module_index: 19, name: L1_Mu6_HTT250er
         15, -- module_index: 20, name: L1_SingleMu12_DQ_EMTF
         32, -- module_index: 21, name: L1_SingleMu16er1p5
         21, -- module_index: 22, name: L1_SingleMu22_OMTF
         28, -- module_index: 23, name: L1_SingleMu9er1p5
        224, -- module_index: 24, name: L1_TripleEG_16_12_8_er2p5
        207, -- module_index: 25, name: L1_DoubleEG_22_10_er2p5
        214, -- module_index: 26, name: L1_DoubleEG_LooseIso22_12_er2p5
        342, -- module_index: 27, name: L1_DoubleJet120er2p5
        188, -- module_index: 28, name: L1_SingleIsoEG28_FWD2p5
        238, -- module_index: 29, name: L1_LooseIsoEG24er2p1_HTT100er
        239, -- module_index: 30, name: L1_LooseIsoEG26er2p1_HTT100er
        241, -- module_index: 31, name: L1_LooseIsoEG30er2p1_HTT100er
        179, -- module_index: 32, name: L1_SingleLooseIsoEG28er2p1
        240, -- module_index: 33, name: L1_LooseIsoEG28er2p1_HTT100er
        186, -- module_index: 34, name: L1_SingleIsoEG26er2p1
        192, -- module_index: 35, name: L1_SingleIsoEG30er2p5
        331, -- module_index: 36, name: L1_SingleJet12erHE
        316, -- module_index: 37, name: L1_SingleJet35er2p5
        175, -- module_index: 38, name: L1_SingleLooseIsoEG26er2p5
        271, -- module_index: 39, name: L1_SingleTau130er2p1
    others => 0
);

-- ========================================================