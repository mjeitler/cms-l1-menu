-- ========================================================
-- from VHDL producer:

-- Module ID: 0

-- Name of L1 Trigger Menu:
-- L1Menu_Collisions2017_dev_r5

-- Unique ID of L1 Trigger Menu:
-- a9c22674-c07e-4484-be32-d1f0726031c7

-- Unique ID of firmware implementation:
-- 38c2787b-f3a1-48e6-b3f8-b7625293f15a

-- Scale set:
-- scales_2017_01_12

-- VHDL producer version
-- v1.0.0

-- HB 2016-09-16: constants for algo_mapping_rop.
type global_index_array is array (0 to NR_ALGOS-1) of integer;
constant global_index: global_index_array := (
        375, -- module_index: 0, name: L1_TripleMu_5_0_0_DoubleMu_5_0_OS_Mass_Max17
         30, -- module_index: 1, name: L1_TripleMu_5_0_0
        415, -- module_index: 2, name: L1_QuadJet36er3p0_Tau52
        151, -- module_index: 3, name: L1_QuadJet50er3p0
        305, -- module_index: 4, name: L1_IsoEG22er2p1_IsoTau26er2p1_dEta_Min0p2
        428, -- module_index: 5, name: L1_Mu3_JetC16_dEta_Max0p4_dPhi_Max0p4
        370, -- module_index: 6, name: L1_DoubleMu0er1p5_SQ_OS_dR_Max1p4
        416, -- module_index: 7, name: L1_ETM75_Jet60_dPhi_Min0p4
        148, -- module_index: 8, name: L1_TripleJet_88_72_56_VBF
        306, -- module_index: 9, name: L1_Mu16er2p1_Tau20er2p1
        307, -- module_index: 10, name: L1_Mu16er2p1_Tau24er2p1
        308, -- module_index: 11, name: L1_Mu18er2p1_Tau20er2p1
         14, -- module_index: 12, name: L1_SingleMu16er2p1
        310, -- module_index: 13, name: L1_Mu18er2p1_IsoTau26er2p1
         15, -- module_index: 14, name: L1_SingleMu18er2p1
        309, -- module_index: 15, name: L1_Mu18er2p1_Tau24er2p1
         16, -- module_index: 16, name: L1_SingleMu20er2p1
        311, -- module_index: 17, name: L1_Mu20er2p1_IsoTau26er2p1
         90, -- module_index: 18, name: L1_DoubleEG_25_14
        108, -- module_index: 19, name: L1_DoubleIsoTau32er2p1
        113, -- module_index: 20, name: L1_DoubleIsoTau38er2p1
        141, -- module_index: 21, name: L1_DoubleJet50er3p0
         27, -- module_index: 22, name: L1_TripleMu0
         32, -- module_index: 23, name: L1_TripleMu_5_5_3
         24, -- module_index: 24, name: L1_DoubleMu_13_6
         44, -- module_index: 25, name: L1_SingleEG24
         48, -- module_index: 26, name: L1_SingleEG32
         51, -- module_index: 27, name: L1_SingleEG38
         68, -- module_index: 28, name: L1_SingleIsoEG18er2p1
         71, -- module_index: 29, name: L1_SingleIsoEG24er2p1
         63, -- module_index: 30, name: L1_SingleIsoEG30
         76, -- module_index: 31, name: L1_SingleIsoEG34er2p1
        126, -- module_index: 32, name: L1_SingleJet140
        121, -- module_index: 33, name: L1_SingleJet20
        101, -- module_index: 34, name: L1_SingleTau80er2p1
         11, -- module_index: 35, name: L1_SingleMu25
        194, -- module_index: 36, name: L1_ETM120
        185, -- module_index: 37, name: L1_ETM75
        171, -- module_index: 38, name: L1_HTT380er
    others => 0
);

-- ========================================================