-- ========================================================
-- from VHDL producer:

-- Module ID: 3

-- Name of L1 Trigger Menu:
-- L1Menu_Collisions2018_v1_0_0

-- Unique ID of L1 Trigger Menu:
-- 409fce06-5701-4b18-9364-39736bfcaf88

-- Unique ID of firmware implementation:
-- 324ed470-bdf0-4315-a64f-da3b4bc3343c

-- Scale set:
-- scales_2017_05_23

-- VHDL producer version
-- v2.3.0

-- HB 2016-09-16: constants for algo_mapping_rop.
type global_index_array is array (0 to NR_ALGOS-1) of integer;
constant global_index: global_index_array := (
        491, -- module_index: 0, name: L1_BPTX_BeamGas_B1_VME
        484, -- module_index: 1, name: L1_BPTX_OR_Ref4_VME
        500, -- module_index: 2, name: L1_HCAL_LaserMon_Trig
        504, -- module_index: 3, name: L1_TOTEM_2
        416, -- module_index: 4, name: L1_ETM120
        411, -- module_index: 5, name: L1_ETT1600
        401, -- module_index: 6, name: L1_HTT255er
        165, -- module_index: 7, name: L1_SingleEG15er2p5
        169, -- module_index: 8, name: L1_SingleEG38er2p5
        173, -- module_index: 9, name: L1_SingleEG50
        183, -- module_index: 10, name: L1_SingleIsoEG24er2p1
        190, -- module_index: 11, name: L1_SingleIsoEG28er1p5
        194, -- module_index: 12, name: L1_SingleIsoEG32er2p1
        319, -- module_index: 13, name: L1_SingleJet120er2p5
        322, -- module_index: 14, name: L1_SingleJet180er2p5
        310, -- module_index: 15, name: L1_SingleJet60
        180, -- module_index: 16, name: L1_SingleLooseIsoEG28er1p5
        238, -- module_index: 17, name: L1_LooseIsoEG24er2p1_HTT100er
        241, -- module_index: 18, name: L1_LooseIsoEG30er2p1_HTT100er
        239, -- module_index: 19, name: L1_LooseIsoEG26er2p1_HTT100er
        240, -- module_index: 20, name: L1_LooseIsoEG28er2p1_HTT100er
        215, -- module_index: 21, name: L1_DoubleEG_LooseIso25_12_er2p5
        341, -- module_index: 22, name: L1_DoubleJet100er2p5
        218, -- module_index: 23, name: L1_DoubleLooseIsoEG24er2p1
        325, -- module_index: 24, name: L1_SingleJet60_FWD3p0
        225, -- module_index: 25, name: L1_TripleEG_16_15_8_er2p5
          5, -- module_index: 26, name: L1_SingleMu0_DQ
         13, -- module_index: 27, name: L1_SingleMu12_DQ_BMTF
         31, -- module_index: 28, name: L1_SingleMu14er1p5
         33, -- module_index: 29, name: L1_SingleMu18er1p5
         21, -- module_index: 30, name: L1_SingleMu22_OMTF
         25, -- module_index: 31, name: L1_SingleMu6er1p5
         26, -- module_index: 32, name: L1_SingleMu7er1p5
          0, -- module_index: 33, name: L1_SingleMuCosmics
        281, -- module_index: 34, name: L1_Mu18er2p1_Tau24er2p1
        282, -- module_index: 35, name: L1_Mu18er2p1_Tau26er2p1
         40, -- module_index: 36, name: L1_DoubleMu0
         42, -- module_index: 37, name: L1_DoubleMu0_SQ_OS
         56, -- module_index: 38, name: L1_DoubleMu0er1p5_SQ_OS
         51, -- module_index: 39, name: L1_DoubleMu18er2p1
         62, -- module_index: 40, name: L1_DoubleMu4p5_SQ_OS
         44, -- module_index: 41, name: L1_DoubleMu9_SQ
         47, -- module_index: 42, name: L1_DoubleMu_15_5_SQ
         49, -- module_index: 43, name: L1_DoubleMu_15_7_SQ
         72, -- module_index: 44, name: L1_TripleMu0
         73, -- module_index: 45, name: L1_TripleMu0_SQ
         75, -- module_index: 46, name: L1_TripleMu3_SQ
         78, -- module_index: 47, name: L1_TripleMu_5_3_3
         79, -- module_index: 48, name: L1_TripleMu_5_3_3_SQ
         77, -- module_index: 49, name: L1_TripleMu_5_3p5_2p5
         83, -- module_index: 50, name: L1_TripleMu_5_3p5_2p5_DoubleMu_5_2p5_OS_Mass_5to17
         84, -- module_index: 51, name: L1_TripleMu_5_4_2p5_DoubleMu_5_2p5_OS_Mass_5to17
         58, -- module_index: 52, name: L1_DoubleMu0er1p5_SQ_OS_dR_Max1p4
         61, -- module_index: 53, name: L1_DoubleMu4_SQ_OS_dR_Max1p2
         50, -- module_index: 54, name: L1_DoubleMu_15_7_Mass_Min1
        356, -- module_index: 55, name: L1_DoubleJet_100_30_DoubleJet30_Mass_Min620
        355, -- module_index: 56, name: L1_DoubleJet_90_30_DoubleJet30_Mass_Min620
        349, -- module_index: 57, name: L1_DoubleJet30er2p5_Mass_Min200_dEta_Max1p5
        257, -- module_index: 58, name: L1_LooseIsoEG22er2p1_IsoTau26er2p1_dR_Min0p3
        236, -- module_index: 59, name: L1_LooseIsoEG30er2p1_Jet34er2p5_dR_Min0p3
        121, -- module_index: 60, name: L1_Mu3_Jet16er2p5_dR_Max0p4
        136, -- module_index: 61, name: L1_Mu12er2p3_Jet40er2p1_dR_Max0p4_DoubleJet40er2p1_dEta_Max1p6
    others => 0
);

-- ========================================================