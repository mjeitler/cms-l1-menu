-- Description:
-- Mapping of algo indexes for ROP

-- ========================================================
-- from VHDL producer:
      
-- Unique ID of L1 Trigger Menu:
-- X"f2fd248d6be8532680fb89a002087e9e"
    
-- Name of L1 Trigger Menu:
-- L1Menu_Collisions2015_25nsStage1_v7_uGT_v4
    
-- Scale set:
-- CMS-IN-2013/XXX
    
-- VHDL producer version
-- v0.0.1

-- ========================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

use work.gtl_pkg.ALL;
use work.gt_mp7_core_pkg.all;

entity algo_mapping_rop is
    port(
        lhc_clk : in std_logic;
        algo_before_prescaler : in std_logic_vector(NR_ALGOS-1 downto 0);
        algo_after_prescaler : in std_logic_vector(NR_ALGOS-1 downto 0);
        algo_after_finor_mask : in std_logic_vector(NR_ALGOS-1 downto 0);
        algo_before_prescaler_rop : out std_logic_vector(MAX_NR_ALGOS-1 downto 0);
        algo_after_prescaler_rop : out std_logic_vector(MAX_NR_ALGOS-1 downto 0);
        algo_after_finor_mask_rop : out std_logic_vector(MAX_NR_ALGOS-1 downto 0)
    );
end algo_mapping_rop;

architecture rtl of algo_mapping_rop is
    signal a_b_p: std_logic_vector(NR_ALGOS-1 downto 0);
    signal a_a_p: std_logic_vector(NR_ALGOS-1 downto 0);
    signal a_a_f: std_logic_vector(NR_ALGOS-1 downto 0);
    signal algo_before_prescaler_rop_int: std_logic_vector(MAX_NR_ALGOS-1 downto 0);
    signal algo_after_prescaler_rop_int: std_logic_vector(MAX_NR_ALGOS-1 downto 0);
    signal algo_after_finor_mask_rop_int: std_logic_vector(MAX_NR_ALGOS-1 downto 0);
begin

a_b_p <= algo_before_prescaler;
a_a_p <= algo_after_prescaler;
a_a_f <= algo_after_finor_mask;

-- ==== Inserted by TME - begin =============================================================================================================

algo_before_prescaler_rop_int <= (
0 => a_b_p(0),
1 => a_b_p(1),
2 => a_b_p(2),
3 => a_b_p(3),
4 => a_b_p(4),
5 => a_b_p(5),
6 => a_b_p(6),
7 => a_b_p(7),
8 => a_b_p(8),
9 => a_b_p(9),
10 => a_b_p(10),
11 => a_b_p(11),
12 => a_b_p(12),
13 => a_b_p(13),
14 => a_b_p(14),
15 => a_b_p(15),
16 => a_b_p(16),
17 => a_b_p(17),
18 => a_b_p(18),
19 => a_b_p(19),
20 => a_b_p(20),
21 => a_b_p(21),
22 => a_b_p(22),
23 => a_b_p(23),
24 => a_b_p(24),
25 => a_b_p(25),
26 => a_b_p(26),
27 => a_b_p(27),
28 => a_b_p(28),
29 => a_b_p(29),
30 => a_b_p(30),
31 => a_b_p(31),
32 => a_b_p(32),
33 => a_b_p(33),
34 => a_b_p(34),
35 => a_b_p(35),
36 => a_b_p(36),
37 => a_b_p(37),
38 => a_b_p(38),
39 => a_b_p(39),
40 => a_b_p(40),
41 => a_b_p(41),
42 => a_b_p(42),
43 => a_b_p(43),
44 => a_b_p(44),
45 => a_b_p(45),
46 => a_b_p(46),
47 => a_b_p(47),
48 => a_b_p(48),
49 => a_b_p(49),
50 => a_b_p(50),
51 => a_b_p(51),
52 => a_b_p(52),
53 => a_b_p(53),
54 => a_b_p(54),
55 => a_b_p(55),
56 => a_b_p(56),
57 => a_b_p(57),
58 => a_b_p(58),
59 => a_b_p(59),
60 => a_b_p(60),
61 => a_b_p(61),
62 => a_b_p(62),
63 => a_b_p(63),
64 => a_b_p(64),
65 => a_b_p(65),
66 => a_b_p(66),
67 => a_b_p(67),
68 => a_b_p(68),
69 => a_b_p(69),
70 => a_b_p(70),
71 => a_b_p(71),
72 => a_b_p(72),
73 => a_b_p(73),
74 => a_b_p(74),
75 => a_b_p(75),
76 => a_b_p(76),
77 => a_b_p(77),
78 => a_b_p(78),
79 => a_b_p(79),
80 => a_b_p(80),
81 => a_b_p(81),
82 => a_b_p(82),
83 => a_b_p(83),
84 => a_b_p(84),
85 => a_b_p(85),
86 => a_b_p(86),
87 => a_b_p(87),
88 => a_b_p(88),
89 => a_b_p(89),
90 => a_b_p(90),
91 => a_b_p(91),
92 => a_b_p(92),
93 => a_b_p(93),
94 => a_b_p(94),
95 => a_b_p(95),
96 => a_b_p(96),
97 => a_b_p(97),
98 => a_b_p(98),
99 => a_b_p(99),
100 => a_b_p(100),
101 => a_b_p(101),
102 => a_b_p(102),
103 => a_b_p(103),
104 => a_b_p(104),
105 => a_b_p(105),
106 => a_b_p(106),
107 => a_b_p(107),
108 => a_b_p(108),
109 => a_b_p(109),
110 => a_b_p(110),
111 => a_b_p(111),
112 => a_b_p(112),
113 => a_b_p(113),
114 => a_b_p(114),
115 => a_b_p(115),
116 => a_b_p(116),
117 => a_b_p(117),
118 => a_b_p(118),
119 => a_b_p(119),
120 => a_b_p(120),
121 => a_b_p(121),
122 => a_b_p(122),
123 => a_b_p(123),
124 => a_b_p(124),
125 => a_b_p(125),
126 => a_b_p(126),
127 => a_b_p(127),
128 => a_b_p(128),
129 => a_b_p(129),
130 => a_b_p(130),
131 => a_b_p(131),
132 => a_b_p(132),
133 => a_b_p(133),
134 => a_b_p(134),
135 => a_b_p(135),
136 => a_b_p(136),
137 => a_b_p(137),
138 => a_b_p(138),
139 => a_b_p(139),
140 => a_b_p(140),
141 => a_b_p(141),
142 => a_b_p(142),
143 => a_b_p(143),
144 => a_b_p(144),
145 => a_b_p(145),
146 => a_b_p(146),
147 => a_b_p(147),
148 => a_b_p(148),
149 => a_b_p(149),
150 => a_b_p(150),
151 => a_b_p(151),
152 => a_b_p(152),
153 => a_b_p(153),
154 => a_b_p(154),
155 => a_b_p(155),
156 => a_b_p(156),
157 => a_b_p(157),
158 => a_b_p(158),
159 => a_b_p(159),
160 => a_b_p(160),
others => '0');

algo_after_prescaler_rop_int <= (
0 => a_a_p(0),
1 => a_a_p(1),
2 => a_a_p(2),
3 => a_a_p(3),
4 => a_a_p(4),
5 => a_a_p(5),
6 => a_a_p(6),
7 => a_a_p(7),
8 => a_a_p(8),
9 => a_a_p(9),
10 => a_a_p(10),
11 => a_a_p(11),
12 => a_a_p(12),
13 => a_a_p(13),
14 => a_a_p(14),
15 => a_a_p(15),
16 => a_a_p(16),
17 => a_a_p(17),
18 => a_a_p(18),
19 => a_a_p(19),
20 => a_a_p(20),
21 => a_a_p(21),
22 => a_a_p(22),
23 => a_a_p(23),
24 => a_a_p(24),
25 => a_a_p(25),
26 => a_a_p(26),
27 => a_a_p(27),
28 => a_a_p(28),
29 => a_a_p(29),
30 => a_a_p(30),
31 => a_a_p(31),
32 => a_a_p(32),
33 => a_a_p(33),
34 => a_a_p(34),
35 => a_a_p(35),
36 => a_a_p(36),
37 => a_a_p(37),
38 => a_a_p(38),
39 => a_a_p(39),
40 => a_a_p(40),
41 => a_a_p(41),
42 => a_a_p(42),
43 => a_a_p(43),
44 => a_a_p(44),
45 => a_a_p(45),
46 => a_a_p(46),
47 => a_a_p(47),
48 => a_a_p(48),
49 => a_a_p(49),
50 => a_a_p(50),
51 => a_a_p(51),
52 => a_a_p(52),
53 => a_a_p(53),
54 => a_a_p(54),
55 => a_a_p(55),
56 => a_a_p(56),
57 => a_a_p(57),
58 => a_a_p(58),
59 => a_a_p(59),
60 => a_a_p(60),
61 => a_a_p(61),
62 => a_a_p(62),
63 => a_a_p(63),
64 => a_a_p(64),
65 => a_a_p(65),
66 => a_a_p(66),
67 => a_a_p(67),
68 => a_a_p(68),
69 => a_a_p(69),
70 => a_a_p(70),
71 => a_a_p(71),
72 => a_a_p(72),
73 => a_a_p(73),
74 => a_a_p(74),
75 => a_a_p(75),
76 => a_a_p(76),
77 => a_a_p(77),
78 => a_a_p(78),
79 => a_a_p(79),
80 => a_a_p(80),
81 => a_a_p(81),
82 => a_a_p(82),
83 => a_a_p(83),
84 => a_a_p(84),
85 => a_a_p(85),
86 => a_a_p(86),
87 => a_a_p(87),
88 => a_a_p(88),
89 => a_a_p(89),
90 => a_a_p(90),
91 => a_a_p(91),
92 => a_a_p(92),
93 => a_a_p(93),
94 => a_a_p(94),
95 => a_a_p(95),
96 => a_a_p(96),
97 => a_a_p(97),
98 => a_a_p(98),
99 => a_a_p(99),
100 => a_a_p(100),
101 => a_a_p(101),
102 => a_a_p(102),
103 => a_a_p(103),
104 => a_a_p(104),
105 => a_a_p(105),
106 => a_a_p(106),
107 => a_a_p(107),
108 => a_a_p(108),
109 => a_a_p(109),
110 => a_a_p(110),
111 => a_a_p(111),
112 => a_a_p(112),
113 => a_a_p(113),
114 => a_a_p(114),
115 => a_a_p(115),
116 => a_a_p(116),
117 => a_a_p(117),
118 => a_a_p(118),
119 => a_a_p(119),
120 => a_a_p(120),
121 => a_a_p(121),
122 => a_a_p(122),
123 => a_a_p(123),
124 => a_a_p(124),
125 => a_a_p(125),
126 => a_a_p(126),
127 => a_a_p(127),
128 => a_a_p(128),
129 => a_a_p(129),
130 => a_a_p(130),
131 => a_a_p(131),
132 => a_a_p(132),
133 => a_a_p(133),
134 => a_a_p(134),
135 => a_a_p(135),
136 => a_a_p(136),
137 => a_a_p(137),
138 => a_a_p(138),
139 => a_a_p(139),
140 => a_a_p(140),
141 => a_a_p(141),
142 => a_a_p(142),
143 => a_a_p(143),
144 => a_a_p(144),
145 => a_a_p(145),
146 => a_a_p(146),
147 => a_a_p(147),
148 => a_a_p(148),
149 => a_a_p(149),
150 => a_a_p(150),
151 => a_a_p(151),
152 => a_a_p(152),
153 => a_a_p(153),
154 => a_a_p(154),
155 => a_a_p(155),
156 => a_a_p(156),
157 => a_a_p(157),
158 => a_a_p(158),
159 => a_a_p(159),
160 => a_a_p(160),
others => '0');

algo_after_finor_mask_rop_int <= (
0 => a_a_f(0),
1 => a_a_f(1),
2 => a_a_f(2),
3 => a_a_f(3),
4 => a_a_f(4),
5 => a_a_f(5),
6 => a_a_f(6),
7 => a_a_f(7),
8 => a_a_f(8),
9 => a_a_f(9),
10 => a_a_f(10),
11 => a_a_f(11),
12 => a_a_f(12),
13 => a_a_f(13),
14 => a_a_f(14),
15 => a_a_f(15),
16 => a_a_f(16),
17 => a_a_f(17),
18 => a_a_f(18),
19 => a_a_f(19),
20 => a_a_f(20),
21 => a_a_f(21),
22 => a_a_f(22),
23 => a_a_f(23),
24 => a_a_f(24),
25 => a_a_f(25),
26 => a_a_f(26),
27 => a_a_f(27),
28 => a_a_f(28),
29 => a_a_f(29),
30 => a_a_f(30),
31 => a_a_f(31),
32 => a_a_f(32),
33 => a_a_f(33),
34 => a_a_f(34),
35 => a_a_f(35),
36 => a_a_f(36),
37 => a_a_f(37),
38 => a_a_f(38),
39 => a_a_f(39),
40 => a_a_f(40),
41 => a_a_f(41),
42 => a_a_f(42),
43 => a_a_f(43),
44 => a_a_f(44),
45 => a_a_f(45),
46 => a_a_f(46),
47 => a_a_f(47),
48 => a_a_f(48),
49 => a_a_f(49),
50 => a_a_f(50),
51 => a_a_f(51),
52 => a_a_f(52),
53 => a_a_f(53),
54 => a_a_f(54),
55 => a_a_f(55),
56 => a_a_f(56),
57 => a_a_f(57),
58 => a_a_f(58),
59 => a_a_f(59),
60 => a_a_f(60),
61 => a_a_f(61),
62 => a_a_f(62),
63 => a_a_f(63),
64 => a_a_f(64),
65 => a_a_f(65),
66 => a_a_f(66),
67 => a_a_f(67),
68 => a_a_f(68),
69 => a_a_f(69),
70 => a_a_f(70),
71 => a_a_f(71),
72 => a_a_f(72),
73 => a_a_f(73),
74 => a_a_f(74),
75 => a_a_f(75),
76 => a_a_f(76),
77 => a_a_f(77),
78 => a_a_f(78),
79 => a_a_f(79),
80 => a_a_f(80),
81 => a_a_f(81),
82 => a_a_f(82),
83 => a_a_f(83),
84 => a_a_f(84),
85 => a_a_f(85),
86 => a_a_f(86),
87 => a_a_f(87),
88 => a_a_f(88),
89 => a_a_f(89),
90 => a_a_f(90),
91 => a_a_f(91),
92 => a_a_f(92),
93 => a_a_f(93),
94 => a_a_f(94),
95 => a_a_f(95),
96 => a_a_f(96),
97 => a_a_f(97),
98 => a_a_f(98),
99 => a_a_f(99),
100 => a_a_f(100),
101 => a_a_f(101),
102 => a_a_f(102),
103 => a_a_f(103),
104 => a_a_f(104),
105 => a_a_f(105),
106 => a_a_f(106),
107 => a_a_f(107),
108 => a_a_f(108),
109 => a_a_f(109),
110 => a_a_f(110),
111 => a_a_f(111),
112 => a_a_f(112),
113 => a_a_f(113),
114 => a_a_f(114),
115 => a_a_f(115),
116 => a_a_f(116),
117 => a_a_f(117),
118 => a_a_f(118),
119 => a_a_f(119),
120 => a_a_f(120),
121 => a_a_f(121),
122 => a_a_f(122),
123 => a_a_f(123),
124 => a_a_f(124),
125 => a_a_f(125),
126 => a_a_f(126),
127 => a_a_f(127),
128 => a_a_f(128),
129 => a_a_f(129),
130 => a_a_f(130),
131 => a_a_f(131),
132 => a_a_f(132),
133 => a_a_f(133),
134 => a_a_f(134),
135 => a_a_f(135),
136 => a_a_f(136),
137 => a_a_f(137),
138 => a_a_f(138),
139 => a_a_f(139),
140 => a_a_f(140),
141 => a_a_f(141),
142 => a_a_f(142),
143 => a_a_f(143),
144 => a_a_f(144),
145 => a_a_f(145),
146 => a_a_f(146),
147 => a_a_f(147),
148 => a_a_f(148),
149 => a_a_f(149),
150 => a_a_f(150),
151 => a_a_f(151),
152 => a_a_f(152),
153 => a_a_f(153),
154 => a_a_f(154),
155 => a_a_f(155),
156 => a_a_f(156),
157 => a_a_f(157),
158 => a_a_f(158),
159 => a_a_f(159),
160 => a_a_f(160),
others => '0');
-- ==== Inserted by TME - end ===============================================================================================================

algo_2_rop_p: process(lhc_clk, algo_before_prescaler_rop_int, algo_after_prescaler_rop_int, algo_after_finor_mask_rop_int)
    begin
    if lhc_clk'event and lhc_clk = '1' then
        algo_before_prescaler_rop <= algo_before_prescaler_rop_int;
        algo_after_prescaler_rop <= algo_after_prescaler_rop_int;
        algo_after_finor_mask_rop <= algo_after_finor_mask_rop_int;
    end if;
end process;

end architecture rtl;