-- ========================================================
-- from VHDL producer:

-- Module ID: 3

-- Name of L1 Trigger Menu:
-- L1Menu_Collisions2017_dev_r5

-- Unique ID of L1 Trigger Menu:
-- a9c22674-c07e-4484-be32-d1f0726031c7

-- Unique ID of firmware implementation:
-- 38c2787b-f3a1-48e6-b3f8-b7625293f15a

-- Scale set:
-- scales_2017_01_12

-- VHDL producer version
-- v1.0.0

-- HB 2016-09-16: constants for algo_mapping_rop.
type global_index_array is array (0 to NR_ALGOS-1) of integer;
constant global_index: global_index_array := (
        371, -- module_index: 0, name: L1_DoubleMu4p5er2p0_SQ_OS_Mass7to18
        423, -- module_index: 1, name: L1_Jet32_Mu0_EG10_dPhi_Jet_Mu_Max0p4_dPhi_Mu_EG_Min1p0
        422, -- module_index: 2, name: L1_Jet32_DoubleMu_10_0_dPhi_Jet_Mu0_Max0p4_dPhi_Mu_Mu_Min1p0
        303, -- module_index: 3, name: L1_IsoEG18er2p1_IsoTau24er2p1_dEta_Min0p2
        253, -- module_index: 4, name: L1_IsoEG30er2p1_Jet34er3p0_dR_Min0p3
        377, -- module_index: 5, name: L1_DoubleMu0er1p4_SQ_OS_dR_Max1p4
        426, -- module_index: 6, name: L1_DoubleMu_10_0_dEta_Max1p8
        376, -- module_index: 7, name: L1_DoubleMu4_OS_EG12
        380, -- module_index: 8, name: L1_DoubleMu5_OS_EG12
         92, -- module_index: 9, name: L1_TripleEG_18_17_8
         84, -- module_index: 10, name: L1_DoubleEG_22_12
         88, -- module_index: 11, name: L1_DoubleEG_25_12
        106, -- module_index: 12, name: L1_DoubleIsoTau28er2p1
        111, -- module_index: 13, name: L1_DoubleIsoTau35er2p1
        146, -- module_index: 14, name: L1_DoubleJet120er3p0
        105, -- module_index: 15, name: L1_DoubleTau70er2p1
         31, -- module_index: 16, name: L1_TripleMu_5_3_3
         23, -- module_index: 17, name: L1_DoubleMu_12_8
         43, -- module_index: 18, name: L1_SingleEG18
         47, -- module_index: 19, name: L1_SingleEG30
         55, -- module_index: 20, name: L1_SingleEG36er2p1
         40, -- module_index: 21, name: L1_SingleEG5
         60, -- module_index: 22, name: L1_SingleIsoEG24
         73, -- module_index: 23, name: L1_SingleIsoEG28er2p1
         65, -- module_index: 24, name: L1_SingleIsoEG34
        125, -- module_index: 25, name: L1_SingleJet120
        130, -- module_index: 26, name: L1_SingleJet180
        100, -- module_index: 27, name: L1_SingleTau20
         17, -- module_index: 28, name: L1_SingleMu22er2p1
        192, -- module_index: 29, name: L1_ETM110
        195, -- module_index: 30, name: L1_ETM150
        206, -- module_index: 31, name: L1_ETMHF150
        172, -- module_index: 32, name: L1_HTT400er
    others => 0
);

-- ========================================================