-- ========================================================
-- from VHDL producer:

-- Module ID: 5

-- Name of L1 Trigger Menu:
-- L1Menu_Collisions2017_dev

-- Unique ID of L1 Trigger Menu:
-- ff279b6e-899e-468b-9704-5fa64b5c005d

-- Unique ID of firmware implementation:
-- 8a4c21f6-5307-4a58-800b-1a1b4e9802a7

-- Scale set:
-- scales_2017_01_12

-- VHDL producer version
-- v1.0.0

-- HB 2016-09-16: constants for algo_mapping_rop.
type global_index_array is array (0 to NR_ALGOS-1) of integer;
constant global_index: global_index_array := (
        374, -- module_index: 0, name: L1_DoubleMu_20_2_SQ_Mass_Max20
        277, -- module_index: 1, name: L1_Mu12er2p3_Jet40er2p3_dR_Max0p4_DoubleJet40er2p3_dEta_Max1p6
        275, -- module_index: 2, name: L1_DoubleJet100er2p3_dEta_Max1p6
        250, -- module_index: 3, name: L1_IsoEG24er2p1_Jet26er3p0_dR_Min0p3
        429, -- module_index: 4, name: L1_Mu3_JetC60_dEta_Max0p4_dPhi_Max0p4
        215, -- module_index: 5, name: L1_CDC_3_TOP_DPHI2p618_3p665
        218, -- module_index: 6, name: L1_CDC_3_er1p6_TOP120_DPHI2p618_3p665
        226, -- module_index: 7, name: L1_CDC_SingleMu_3_er1p6_TOP120_DPHI2p618_3p665
        377, -- module_index: 8, name: L1_DoubleMu0er1p4_SQ_OS_dR_Max1p4
        289, -- module_index: 9, name: L1_ETM100_Jet60_dPhi_Min0p4
        287, -- module_index: 10, name: L1_ETM80_Jet60_dPhi_Min0p4
        149, -- module_index: 11, name: L1_TripleJet_92_76_64_VBF
         80, -- module_index: 12, name: L1_DoubleEG_15_10
         83, -- module_index: 13, name: L1_DoubleEG_22_10
         88, -- module_index: 14, name: L1_DoubleEG_25_12
        106, -- module_index: 15, name: L1_DoubleIsoTau28er2p1
        111, -- module_index: 16, name: L1_DoubleIsoTau35er2p1
        146, -- module_index: 17, name: L1_DoubleJet120er3p0
        105, -- module_index: 18, name: L1_DoubleTau70er2p1
         32, -- module_index: 19, name: L1_TripleMu_5_5_3
         26, -- module_index: 20, name: L1_DoubleMu_15_7
         46, -- module_index: 21, name: L1_SingleEG28
         50, -- module_index: 22, name: L1_SingleEG36
         53, -- module_index: 23, name: L1_SingleEG45
         70, -- module_index: 24, name: L1_SingleIsoEG22er2p1
         62, -- module_index: 25, name: L1_SingleIsoEG28
         75, -- module_index: 26, name: L1_SingleIsoEG32er2p1
         67, -- module_index: 27, name: L1_SingleIsoEG38
        128, -- module_index: 28, name: L1_SingleJet160
        102, -- module_index: 29, name: L1_SingleTau100er2p1
          7, -- module_index: 30, name: L1_SingleMu16
         12, -- module_index: 31, name: L1_SingleMu30
        193, -- module_index: 32, name: L1_ETM115
        185, -- module_index: 33, name: L1_ETM75
        170, -- module_index: 34, name: L1_HTT340er
    others => 0
);

-- ========================================================