-- ========================================================
-- from VHDL producer:

-- Module ID: 0

-- Name of L1 Trigger Menu:
-- L1Menu_Collisions2017_dev

-- Unique ID of L1 Trigger Menu:
-- ff279b6e-899e-468b-9704-5fa64b5c005d

-- Unique ID of firmware implementation:
-- 8a4c21f6-5307-4a58-800b-1a1b4e9802a7

-- Scale set:
-- scales_2017_01_12

-- VHDL producer version
-- v1.0.0

-- HB 2016-09-16: constants for algo_mapping_rop.
type global_index_array is array (0 to NR_ALGOS-1) of integer;
constant global_index: global_index_array := (
        375, -- module_index: 0, name: L1_TripleMu_5_0_0_DoubleMu_5_0_OS_Mass_Max17
         30, -- module_index: 1, name: L1_TripleMu_5_0_0
        415, -- module_index: 2, name: L1_QuadJet36er3p0_Tau52
        151, -- module_index: 3, name: L1_QuadJet50er3p0
        305, -- module_index: 4, name: L1_IsoEG22er2p1_IsoTau26er2p1_dEta_Min0p2
        428, -- module_index: 5, name: L1_Mu3_JetC16_dEta_Max0p4_dPhi_Max0p4
        216, -- module_index: 6, name: L1_CDC_3_TOP120_DPHI2p618_3p665
        222, -- module_index: 7, name: L1_CDC_3_er1p6_TOP120_DPHI2p094_4p189
        227, -- module_index: 8, name: L1_CDC_SingleMu_3_er1p2_TOP120_DPHI2p618_3p665
        229, -- module_index: 9, name: L1_CDCp1_3_er2p1_TOP120_DPHI2p618_3p665
        426, -- module_index: 10, name: L1_DoubleMu_10_0_dEta_Max1p8
        376, -- module_index: 11, name: L1_DoubleMu4_OS_EG12
        380, -- module_index: 12, name: L1_DoubleMu5_OS_EG12
        306, -- module_index: 13, name: L1_Mu16er2p1_Tau20er2p1
        310, -- module_index: 14, name: L1_Mu18er2p1_IsoTau26er2p1
        307, -- module_index: 15, name: L1_Mu16er2p1_Tau24er2p1
         16, -- module_index: 16, name: L1_SingleMu20er2p1
        311, -- module_index: 17, name: L1_Mu20er2p1_IsoTau26er2p1
        308, -- module_index: 18, name: L1_Mu18er2p1_Tau20er2p1
         15, -- module_index: 19, name: L1_SingleMu18er2p1
        309, -- module_index: 20, name: L1_Mu18er2p1_Tau24er2p1
         14, -- module_index: 21, name: L1_SingleMu16er2p1
         85, -- module_index: 22, name: L1_DoubleEG_22_15
         90, -- module_index: 23, name: L1_DoubleEG_25_14
        108, -- module_index: 24, name: L1_DoubleIsoTau32er2p1
        113, -- module_index: 25, name: L1_DoubleIsoTau38er2p1
        141, -- module_index: 26, name: L1_DoubleJet50er3p0
         27, -- module_index: 27, name: L1_TripleMu0
        381, -- module_index: 28, name: L1_DoubleMu6_SQ_OS
         24, -- module_index: 29, name: L1_DoubleMu_13_6
         44, -- module_index: 30, name: L1_SingleEG24
         48, -- module_index: 31, name: L1_SingleEG32
         51, -- module_index: 32, name: L1_SingleEG38
         68, -- module_index: 33, name: L1_SingleIsoEG18er2p1
         71, -- module_index: 34, name: L1_SingleIsoEG24er2p1
         63, -- module_index: 35, name: L1_SingleIsoEG30
         76, -- module_index: 36, name: L1_SingleIsoEG34er2p1
        126, -- module_index: 37, name: L1_SingleJet140
        121, -- module_index: 38, name: L1_SingleJet20
          5, -- module_index: 39, name: L1_SingleMu10_LowQ
         11, -- module_index: 40, name: L1_SingleMu25
        191, -- module_index: 41, name: L1_ETM105
        195, -- module_index: 42, name: L1_ETM150
        160, -- module_index: 43, name: L1_HTT120er
        172, -- module_index: 44, name: L1_HTT400er
    others => 0
);

-- ========================================================