-- ========================================================
-- from VHDL producer:

-- Module ID: 0

-- Name of L1 Trigger Menu:
-- L1Menu_CollisionsHeavyIons2018_v3

-- Unique ID of L1 Trigger Menu:
-- bb9a82eb-17df-4991-b806-4028ee613a4c

-- Unique ID of firmware implementation:
-- 721d74e7-03e3-48ab-938d-1e8242e7c1dd

-- Scale set:
-- scales_2018_08_07

-- VHDL producer version
-- v2.5.0

-- HB 2016-09-16: constants for algo_mapping_rop.
type global_index_array is array (0 to NR_ALGOS-1) of integer;
constant global_index: global_index_array := (
        296, -- module_index: 0, name: L1_DoubleMuOpen_MaxDr2p0_BptxAND
          9, -- module_index: 1, name: L1_AlwaysTrue
          1, -- module_index: 2, name: L1_ZeroBias_copy
          0, -- module_index: 3, name: L1_ZeroBias
    others => 0
);

-- ========================================================