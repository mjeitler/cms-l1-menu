-- ========================================================
-- from VHDL producer:

-- Module ID: 1

-- Name of L1 Trigger Menu:
-- L1Menu_Collisions2017_dev

-- Unique ID of L1 Trigger Menu:
-- a062fa36-6b9d-4302-9842-2e606a849e32

-- Unique ID of firmware implementation:
-- d2bef55e-4757-4a07-8032-f42a7daea756

-- Scale set:
-- scales_2017_01_12

-- VHDL producer version
-- v1.0.0

-- HB 2016-09-16: constants for algo_mapping_rop.
type global_index_array is array (0 to NR_ALGOS-1) of integer;
constant global_index: global_index_array := (
        359, -- module_index: 0, name: L1_TripleMu_5_3_0_DoubleMu_5_3_OS_Mass_Max17
        281, -- module_index: 1, name: L1_Mu10er2p3_Jet32er2p3_dR_Max0p4_DoubleJet32er2p3_dEta_Max1p6
        434, -- module_index: 2, name: L1_QuadJet36er3p0_Tau52
        151, -- module_index: 3, name: L1_QuadJet50er3p0
        295, -- module_index: 4, name: L1_IsoEG18er2p1_IsoTau24er2p1_dEta_Min0p2
        261, -- module_index: 5, name: L1_IsoEG26er2p1_Jet30er3p0_dR_Min0p3
        404, -- module_index: 6, name: L1_Mu3_JetC60_dEta_Max0p4_dPhi_Max0p4
        350, -- module_index: 7, name: L1_DoubleMu0er1p5_SQ_OS_dR_Max1p4
        286, -- module_index: 8, name: L1_ETM100cer_Jet60_dPhi_Min0p4
        435, -- module_index: 9, name: L1_ETM75cer_Jet60_dPhi_Min0p4
        147, -- module_index: 10, name: L1_TripleJet_84_68_48_VBF
         33, -- module_index: 11, name: L1_QuadMu0
         91, -- module_index: 12, name: L1_TripleEG_14_10_8
        287, -- module_index: 13, name: L1_DoubleJet60er3p0_ETM80cer
        186, -- module_index: 14, name: L1_ETM80cer
         81, -- module_index: 15, name: L1_DoubleEG_18_17
         84, -- module_index: 16, name: L1_DoubleEG_22_12
         87, -- module_index: 17, name: L1_DoubleEG_24_17
         90, -- module_index: 18, name: L1_DoubleEG_25_14
        105, -- module_index: 19, name: L1_DoubleIsoTau28er2p1
        108, -- module_index: 20, name: L1_DoubleIsoTau33er2p1
        112, -- module_index: 21, name: L1_DoubleIsoTau38er2p1
        140, -- module_index: 22, name: L1_DoubleJet40er3p0
        104, -- module_index: 23, name: L1_DoubleTau70er2p1
         29, -- module_index: 24, name: L1_TripleMu_4_4_4
         21, -- module_index: 25, name: L1_DoubleMu_11_4
         24, -- module_index: 26, name: L1_DoubleMu_13_6
        414, -- module_index: 27, name: L1_Mu8_HTT150er
         45, -- module_index: 28, name: L1_SingleEG26
         48, -- module_index: 29, name: L1_SingleEG32
         50, -- module_index: 30, name: L1_SingleEG36
         56, -- module_index: 31, name: L1_SingleEG38er2p1
         40, -- module_index: 32, name: L1_SingleEG5
         59, -- module_index: 33, name: L1_SingleIsoEG22
         71, -- module_index: 34, name: L1_SingleIsoEG24er2p1
         73, -- module_index: 35, name: L1_SingleIsoEG28er2p1
         75, -- module_index: 36, name: L1_SingleIsoEG32er2p1
         77, -- module_index: 37, name: L1_SingleIsoEG36er2p1
        127, -- module_index: 38, name: L1_SingleJet150
        130, -- module_index: 39, name: L1_SingleJet180
        101, -- module_index: 40, name: L1_SingleTau100er2p1
          6, -- module_index: 41, name: L1_SingleMu11_LowQ
         17, -- module_index: 42, name: L1_SingleMu22er2p1
          0, -- module_index: 43, name: L1_SingleMuCosmics
        185, -- module_index: 44, name: L1_ETM75cer
        206, -- module_index: 45, name: L1_ETMHF150c
        170, -- module_index: 46, name: L1_HTT340er
        174, -- module_index: 47, name: L1_HTT500er
    others => 0
);

-- ========================================================