-- ========================================================
-- from VHDL producer:

-- Module ID: 3

-- Name of L1 Trigger Menu:
-- L1Menu_Collisions2017_dev

-- Unique ID of L1 Trigger Menu:
-- ff279b6e-899e-468b-9704-5fa64b5c005d

-- Unique ID of firmware implementation:
-- 8a4c21f6-5307-4a58-800b-1a1b4e9802a7

-- Scale set:
-- scales_2017_01_12

-- VHDL producer version
-- v1.0.0

-- HB 2016-09-16: constants for algo_mapping_rop.
type global_index_array is array (0 to NR_ALGOS-1) of integer;
constant global_index: global_index_array := (
        371, -- module_index: 0, name: L1_DoubleMu4p5er2p0_SQ_OS_Mass7to18
        423, -- module_index: 1, name: L1_Jet32_Mu0_EG10_dPhi_Jet_Mu_Max0p4_dPhi_Mu_EG_Min1p0
        422, -- module_index: 2, name: L1_Jet32_DoubleMu_10_0_dPhi_Jet_Mu0_Max0p4_dPhi_Mu_Mu_Min1p0
        303, -- module_index: 3, name: L1_IsoEG18er2p1_IsoTau24er2p1_dEta_Min0p2
        253, -- module_index: 4, name: L1_IsoEG30er2p1_Jet34er3p0_dR_Min0p3
        232, -- module_index: 5, name: L1_CDC_3_TOP120_DPHI1p570_4p711
        223, -- module_index: 6, name: L1_CDC_3_er1p2_TOP120_DPHI2p094_4p189
        221, -- module_index: 7, name: L1_CDC_3_er2p1_TOP120_DPHI2p094_4p189
        228, -- module_index: 8, name: L1_CDCp1_3_TOP120_DPHI2p618_3p665
        370, -- module_index: 9, name: L1_DoubleMu0er1p5_SQ_OS_dR_Max1p4
        416, -- module_index: 10, name: L1_ETM75_Jet60_dPhi_Min0p4
        148, -- module_index: 11, name: L1_TripleJet_88_72_56_VBF
        297, -- module_index: 12, name: L1_TripleEG_Iso20_10_5
         86, -- module_index: 13, name: L1_DoubleEG_23_10
        295, -- module_index: 14, name: L1_DoubleEG_Iso23_10
        109, -- module_index: 15, name: L1_DoubleIsoTau33er2p1
        144, -- module_index: 16, name: L1_DoubleJet100er3p0
        143, -- module_index: 17, name: L1_DoubleJet80er3p0
         28, -- module_index: 18, name: L1_TripleMu3
         21, -- module_index: 19, name: L1_DoubleMu_11_4
        438, -- module_index: 20, name: L1_Mu10er2p1_ETM30
        439, -- module_index: 21, name: L1_Mu14er2p1_ETM30
        180, -- module_index: 22, name: L1_ETM30
         13, -- module_index: 23, name: L1_SingleMu14er2p1
         49, -- module_index: 24, name: L1_SingleEG34
         56, -- module_index: 25, name: L1_SingleEG38er2p1
         69, -- module_index: 26, name: L1_SingleIsoEG20er2p1
         61, -- module_index: 27, name: L1_SingleIsoEG26
         74, -- module_index: 28, name: L1_SingleIsoEG30er2p1
         66, -- module_index: 29, name: L1_SingleIsoEG36
        127, -- module_index: 30, name: L1_SingleJet150
        131, -- module_index: 31, name: L1_SingleJet200
        101, -- module_index: 32, name: L1_SingleTau80er2p1
          0, -- module_index: 33, name: L1_SingleMuCosmics
        194, -- module_index: 34, name: L1_ETM120
        206, -- module_index: 35, name: L1_ETMHF150
        171, -- module_index: 36, name: L1_HTT380er
    others => 0
);

-- ========================================================